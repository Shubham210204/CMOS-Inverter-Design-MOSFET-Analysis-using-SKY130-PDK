magic
tech sky130A
timestamp 1742055881
<< nwell >>
rect -200 -120 100 200
<< nmos >>
rect -60 -285 -45 -185
<< pmos >>
rect -60 -100 -45 100
<< ndiff >>
rect -105 -225 -60 -185
rect -105 -245 -95 -225
rect -75 -245 -60 -225
rect -105 -285 -60 -245
rect -45 -225 0 -185
rect -45 -245 -30 -225
rect -10 -245 0 -225
rect -45 -285 0 -245
<< pdiff >>
rect -105 10 -60 100
rect -105 -10 -95 10
rect -75 -10 -60 10
rect -105 -100 -60 -10
rect -45 10 0 100
rect -45 -10 -30 10
rect -10 -10 0 10
rect -45 -100 0 -10
<< ndiffc >>
rect -95 -245 -75 -225
rect -30 -245 -10 -225
<< pdiffc >>
rect -95 -10 -75 10
rect -30 -10 -10 10
<< psubdiff >>
rect -105 -330 0 -315
rect -105 -350 -90 -330
rect -70 -350 -35 -330
rect -15 -350 0 -330
rect -105 -365 0 -350
<< nsubdiff >>
rect -105 165 -5 180
rect -105 145 -90 165
rect -70 145 -35 165
rect -15 145 -5 165
rect -105 130 -5 145
<< psubdiffcont >>
rect -90 -350 -70 -330
rect -35 -350 -15 -330
<< nsubdiffcont >>
rect -90 145 -70 165
rect -35 145 -15 165
<< poly >>
rect -60 100 -45 120
rect -60 -125 -45 -100
rect -100 -135 -45 -125
rect -100 -155 -90 -135
rect -70 -155 -45 -135
rect -100 -165 -45 -155
rect -60 -185 -45 -165
rect -60 -305 -45 -285
<< polycont >>
rect -90 -155 -70 -135
<< locali >>
rect -105 165 -5 180
rect -105 145 -90 165
rect -70 145 -35 165
rect -15 145 -5 165
rect -105 130 -5 145
rect -105 10 -65 130
rect -105 -10 -95 10
rect -75 -10 -65 10
rect -105 -100 -65 -10
rect -40 10 0 100
rect -40 -10 -30 10
rect -10 -10 0 10
rect -100 -135 -60 -125
rect -100 -155 -90 -135
rect -70 -155 -60 -135
rect -100 -165 -60 -155
rect -40 -130 0 -10
rect -40 -150 -30 -130
rect -10 -150 0 -130
rect -105 -225 -65 -185
rect -105 -245 -95 -225
rect -75 -245 -65 -225
rect -105 -315 -65 -245
rect -40 -225 0 -150
rect -40 -245 -30 -225
rect -10 -245 0 -225
rect -40 -285 0 -245
rect -105 -330 0 -315
rect -105 -350 -90 -330
rect -70 -350 -35 -330
rect -15 -350 0 -330
rect -105 -365 0 -350
<< viali >>
rect -90 145 -70 165
rect -90 -155 -70 -135
rect -30 -150 -10 -130
rect -90 -350 -70 -330
<< metal1 >>
rect -240 165 140 180
rect -240 145 -90 165
rect -70 145 140 165
rect -240 130 140 145
rect -240 -135 -60 -125
rect -240 -155 -90 -135
rect -70 -155 -60 -135
rect -240 -165 -60 -155
rect -40 -130 140 -120
rect -40 -150 -30 -130
rect -10 -150 140 -130
rect -40 -160 140 -150
rect -240 -330 140 -315
rect -240 -350 -90 -330
rect -70 -350 140 -330
rect -240 -365 140 -350
<< labels >>
rlabel metal1 115 155 115 155 1 vdd
rlabel metal1 115 -345 115 -345 1 gnd
rlabel metal1 140 -160 140 -120 7 output
rlabel metal1 -240 -165 -240 -125 3 input
<< end >>
